library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.all;
use IEEE.NUMERIC_STD.ALL;

entity my_rom_dp_v2 is 
generic(

addr_len: natural := 10;
data_len: natural := 20
);
port(
rom_enable: in std_logic;
address: in std_logic_vector((addr_len -1) downto 0);
data_out: out std_logic_vector((data_len -1) downto 0)
);
end entity;


architecture arch of my_rom_dp_v2 is

type rom_type is array (0 to (2**(addr_len) -1)) of std_logic_vector((data_len -1) downto 0);

constant mem: rom_type := 
	(
	"11111111110000000000",
	
    "11111111010000000110",

    "11111110110000010010",

    "11111110010000100100",

    "11111101110000111100",

    "11111101010001011010",

    "11111100110001111101",

    "11111100010010100111",

    "11111011110011010110",

    "11111011010100001011",

    "11111010110101000110",

    "11111010010110000110",

    "11111001110111001101",

    "11111001011000011001",

    "11111000111001101011",

    "11111000011011000010",

    "11110111111100011111",

    "11110111011110000010",

    "11110110111111101010",

    "11110110100001011000",

    "11110110000011001011",

    "11110101100101000100",

    "11110101000111000011",

    "11110100101001000111",

    "11110100001011010000",

    "11110011101101011111",

    "11110011001111110100",

    "11110010110010001110",

    "11110010010100101101",

    "11110001110111010001",

    "11110001011001111011",

    "11110000111100101011",

    "11110000011111011111",

    "11110000000010011001",

    "11101111100101011000",

    "11101111001000011101",

    "11101110101011100110",

    "11101110001110110101",

    "11101101110010001001",

    "11101101010101100011",

    "11101100111001000001",

    "11101100011100100101",

    "11101100000000001101",

    "11101011100011111011",

    "11101011000111101110",

    "11101010101011100110",

    "11101010001111100011",

    "11101001110011100101",

    "11101001010111101100",

    "11101000111011111000",

    "11101000100000001000",

    "11101000000100011110",

    "11100111101000111001",

    "11100111001101011001",

    "11100110110001111101",

    "11100110010110100111",

    "11100101111011010101",

    "11100101100000001000",

    "11100101000101000000",

    "11100100101001111101",

    "11100100001110111111",

    "11100011110100000101",

    "11100011011001010000",

    "11100010111110100000",

    "11100010100011110101",

    "11100010001001001110",

    "11100001101110101100",

    "11100001010100001111",

    "11100000111001110110",

    "11100000011111100010",

    "11100000000101010010",

    "11011111101011000111",

    "11011111010001000001",

    "11011110110110111111",

    "11011110011101000010",

    "11011110000011001001",

    "11011101101001010101",

    "11011101001111100110",

    "11011100110101111010",

    "11011100011100010100",

    "11011100000010110001",

    "11011011101001010100",

    "11011011001111111010",

    "11011010110110100101",

    "11011010011101010101",

    "11011010000100001000",

    "11011001101011000000",

    "11011001010001111101",

    "11011000111000111110",

    "11011000100000000011",

    "11011000000111001100",

    "11010111101110011010",

    "11010111010101101011",

    "11010110111101000010",

    "11010110100100011100",

    "11010110001011111011",

    "11010101110011011101",

    "11010101011011000100",

    "11010101000010101111",

    "11010100101010011111",

    "11010100010010010010",

    "11010011111010001010",

    "11010011100010000101",

    "11010011001010000101",

    "11010010110010001001",

    "11010010011010010001",

    "11010010000010011101",

    "11010001101010101101",

    "11010001010011000001",

    "11010000111011011001",

    "11010000100011110101",

    "11010000001100010101",

    "11001111110100111001",

    "11001111011101100001",

    "11001111000110001101",

    "11001110101110111101",

    "11001110010111110000",

    "11001110000000101000",

    "11001101101001100011",

    "11001101010010100011",

    "11001100111011100110",

    "11001100100100101101",

    "11001100001101111000",

    "11001011110111000111",

    "11001011100000011001",

    "11001011001001110000",

    "11001010110011001010",

    "11001010011100101000",

    "11001010000110001001",

    "11001001101111101111",

    "11001001011001011000",

    "11001001000011000101",

    "11001000101100110101",

    "11001000010110101001",

    "11001000000000100001",

    "11000111101010011101",

    "11000111010100011100",

    "11000110111110011111",

    "11000110101000100101",

    "11000110010010101111",

    "11000101111100111101",

    "11000101100111001110",

    "11000101010001100011",

    "11000100111011111011",

    "11000100100110010111",

    "11000100010000110111",

    "11000011111011011010",

    "11000011100110000000",

    "11000011010000101010",

    "11000010111011011000",

    "11000010100110001001",

    "11000010010000111101",

    "11000001111011110101",

    "11000001100110110000",

    "11000001010001101111",

    "11000000111100110001",

    "11000000100111110111",

    "11000000010011000000",

    "10111111111110001100",

    "10111111101001011100",

    "10111111010100101111",

    "10111111000000000110",

    "10111110101011011111",

    "10111110010110111101",

    "10111110000010011101",

    "10111101101110000001",

    "10111101011001101000",

    "10111101000101010010",

    "10111100110001000000",

    "10111100011100110001",

    "10111100001000100101",

    "10111011110100011100",

    "10111011100000010111",

    "10111011001100010101",

    "10111010111000010110",

    "10111010100100011010",

    "10111010010000100001",

    "10111001111100101100",

    "10111001101000111010",

    "10111001010101001011",

    "10111001000001011111",

    "10111000101101110110",

    "10111000011010010000",

    "10111000000110101110",

    "10110111110011001110",

    "10110111011111110010",

    "10110111001100011000",

    "10110110111001000010",

    "10110110100101101111",

    "10110110010010011111",

    "10110101111111010010",

    "10110101101100001000",

    "10110101011001000001",

    "10110101000101111101",

    "10110100110010111100",

    "10110100011111111110",

    "10110100001101000011",

    "10110011111010001011",

    "10110011100111010110",

    "10110011010100100100",

    "10110011000001110100",

    "10110010101111001000",

    "10110010011100011111",

    "10110010001001111000",

    "10110001110111010101",

    "10110001100100110100",

    "10110001010010010111",

    "10110000111111111100",

    "10110000101101100100",

    "10110000011011001111",

    "10110000001000111100",

    "10101111110110101101",

    "10101111100100100000",

    "10101111010010010111",

    "10101111000000010000",

    "10101110101110001100",

    "10101110011100001010",

    "10101110001010001100",

    "10101101111000010000",

    "10101101100110010111",

    "10101101010100100001",

    "10101101000010101101",

    "10101100110000111100",

    "10101100011111001110",

    "10101100001101100011",

    "10101011111011111010",

    "10101011101010010100",

    "10101011011000110001",

    "10101011000111010001",

    "10101010110101110011",

    "10101010100100011000",

    "10101010010010111111",

    "10101010000001101001",

    "10101001110000010110",

    "10101001011111000110",

    "10101001001101111000",

    "10101000111100101100",

    "10101000101011100100",

    "10101000011010011110",

    "10101000001001011010",

    "10100111111000011001",

    "10100111100111011011",

    "10100111010110011111",

    "10100111000101100110",

    "10100110110100101111",

    "10100110100011111011",

    "10100110010011001010",

    "10100110000010011011",

    "10100101110001101110",

    "10100101100001000100",

    "10100101010000011101",

    "10100100111111111000",

    "10100100101111010101",

    "10100100011110110101",

    "10100100001110011000",

    "10100011111101111101",

    "10100011101101100100",

    "10100011011101001110",

    "10100011001100111010",

    "10100010111100101001",

    "10100010101100011010",

    "10100010011100001110",

    "10100010001100000100",

    "10100001111011111100",

    "10100001101011110111",

    "10100001011011110100",

    "10100001001011110100",

    "10100000111011110110",

    "10100000101011111010",

    "10100000011100000001",

    "10100000001100001010",

    "10011111111100010110",

    "10011111101100100100",

    "10011111011100110100",

    "10011111001101000110",

    "10011110111101011011",

    "10011110101101110010",

    "10011110011110001011",

    "10011110001110100111",

    "10011101111111000101",

    "10011101101111100101",

    "10011101100000001000",

    "10011101010000101101",

    "10011101000001010100",

    "10011100110001111101",

    "10011100100010101001",

    "10011100010011010110",

    "10011100000100000110",

    "10011011110100111001",

    "10011011100101101101",

    "10011011010110100100",

    "10011011000111011101",

    "10011010111000011000",

    "10011010101001010101",

    "10011010011010010101",

    "10011010001011010111",

    "10011001111100011011",

    "10011001101101100001",

    "10011001011110101001",

    "10011001001111110011",

    "10011001000001000000",

    "10011000110010001110",

    "10011000100011011111",

    "10011000010100110010",

    "10011000000110000111",

    "10010111110111011110",

    "10010111101000111000",

    "10010111011010010011",

    "10010111001011110001",

    "10010110111101010000",

    "10010110101110110010",

    "10010110100000010110",

    "10010110010001111011",

    "10010110000011100011",

    "10010101110101001101",

    "10010101100110111001",

    "10010101011000100111",

    "10010101001010011000",

    "10010100111100001010",

    "10010100101101111110",

    "10010100011111110100",

    "10010100010001101100",

    "10010100000011100110",

    "10010011110101100011",

    "10010011100111100001",

    "10010011011001100001",

    "10010011001011100011",

    "10010010111101101000",

    "10010010101111101110",

    "10010010100001110110",

    "10010010010100000000",

    "10010010000110001100",

    "10010001111000011010",

    "10010001101010101010",

    "10010001011100111100",

    "10010001001111010000",

    "10010001000001100110",

    "10010000110011111110",

    "10010000100110010111",

    "10010000011000110011",

    "10010000001011010000",

    "10001111111101110000",

    "10001111110000010001",

    "10001111100010110100",

    "10001111010101011001",

    "10001111001000000000",

    "10001110111010101001",

    "10001110101101010011",

    "10001110100000000000",

    "10001110010010101110",

    "10001110000101011111",

    "10001101111000010001",

    "10001101101011000101",

    "10001101011101111010",

    "10001101010000110010",

    "10001101000011101011",

    "10001100110110100111",

    "10001100101001100100",

    "10001100011100100011",

    "10001100001111100011",

    "10001100000010100110",

    "10001011110101101010",

    "10001011101000110000",

    "10001011011011111000",

    "10001011001111000010",

    "10001011000010001101",

    "10001010110101011010",

    "10001010101000101001",

    "10001010011011111010",

    "10001010001111001100",

    "10001010000010100001",

    "10001001110101110111",

    "10001001101001001110",

    "10001001011100101000",

    "10001001010000000011",

    "10001001000011100000",

    "10001000110110111110",

    "10001000101010011111",

    "10001000011110000001",

    "10001000010001100100",

    "10001000000101001010",

    "10000111111000110001",

    "10000111101100011010",

    "10000111100000000100",

    "10000111010011110001",

    "10000111000111011110",

    "10000110111011001110",

    "10000110101110111111",

    "10000110100010110010",

    "10000110010110100111",

    "10000110001010011101",

    "10000101111110010101",

    "10000101110010001110",

    "10000101100110001001",

    "10000101011010000110",

    "10000101001110000100",

    "10000101000010000100",

    "10000100110110000110",

    "10000100101010001001",

    "10000100011110001110",

    "10000100010010010100",

    "10000100000110011100",

    "10000011111010100110",

    "10000011101110110001",

    "10000011100010111110",

    "10000011010111001100",

    "10000011001011011100",

    "10000010111111101110",

    "10000010110100000001",

    "10000010101000010110",

    "10000010011100101100",

    "10000010010001000100",

    "10000010000101011101",

    "10000001111001111000",

    "10000001101110010101",

    "10000001100010110011",

    "10000001010111010010",

    "10000001001011110011",

    "10000001000000010110",

    "10000000110100111010",

    "10000000101001100000",

    "10000000011110000111",

    "10000000010010110000",

    "10000000000111011010",

    "11111111111000001100",

    "11111111100001100110",

    "11111111001011000011",

    "11111110110100100100",

    "11111110011110000111",

    "11111110000111101101",

    "11111101110001010111",

    "11111101011011000011",

    "11111101000100110010",

    "11111100101110100100",

    "11111100011000011001",

    "11111100000010010001",

    "11111011101100001100",

    "11111011010110001001",

    "11111011000000001010",

    "11111010101010001101",

    "11111010010100010100",

    "11111001111110011101",

    "11111001101000101001",

    "11111001010010111000",

    "11111000111101001010",

    "11111000100111011110",

    "11111000010001110110",

    "11110111111100010000",

    "11110111100110101101",

    "11110111010001001101",

    "11110110111011110000",

    "11110110100110010101",

    "11110110010000111110",

    "11110101111011101001",

    "11110101100110010110",

    "11110101010001000111",

    "11110100111011111010",

    "11110100100110110000",

    "11110100010001101001",

    "11110011111100100101",

    "11110011100111100011",

    "11110011010010100100",

    "11110010111101101000",

    "11110010101000101110",

    "11110010010011110111",

    "11110001111111000011",

    "11110001101010010001",

    "11110001010101100011",

    "11110001000000110110",

    "11110000101100001101",

    "11110000010111100110",

    "11110000000011000010",

    "11101111101110100000",

    "11101111011010000001",

    "11101111000101100101",

    "11101110110001001011",

    "11101110011100110100",

    "11101110001000011111",

    "11101101110100001101",

    "11101101011111111110",

    "11101101001011110001",

    "11101100110111100111",

    "11101100100011100000",

    "11101100001111011011",

    "11101011111011011000",

    "11101011100111011000",

    "11101011010011011011",

    "11101010111111100000",

    "11101010101011100111",

    "11101010010111110010",

    "11101010000011111110",

    "11101001110000001110",

    "11101001011100011111",

    "11101001001000110011",

    "11101000110101001010",

    "11101000100001100011",

    "11101000001101111111",

    "11100111111010011101",

    "11100111100110111110",

    "11100111010011100001",

    "11100111000000000110",

    "11100110101100101110",

    "11100110011001011000",

    "11100110000110000101",

    "11100101110010110100",

    "11100101011111100110",

    "11100101001100011010",

    "11100100111001010000",

    "11100100100110001001",

    "11100100010011000101",

    "11100100000000000010",

    "11100011101101000010",

    "11100011011010000101",

    "11100011000111001001",

    "11100010110100010000",

    "11100010100001011010",

    "11100010001110100110",

    "11100001111011110100",

    "11100001101001000100",

    "11100001010110010111",

    "11100001000011101100",

    "11100000110001000100",

    "11100000011110011101",

    "11100000001011111010",

    "11011111111001011000",

    "11011111100110111001",

    "11011111010100011100",

    "11011111000010000001",

    "11011110101111101000",

    "11011110011101010010",

    "11011110001010111110",

    "11011101111000101100",

    "11011101100110011101",

    "11011101010100010000",

    "11011101000010000101",

    "11011100101111111100",

    "11011100011101110110",

    "11011100001011110001",

    "11011011111001101111",

    "11011011100111110000",

    "11011011010101110010",

    "11011011000011110111",

    "11011010110001111101",

    "11011010100000000110",

    "11011010001110010010",

    "11011001111100011111",

    "11011001101010101110",

    "11011001011001000000",

    "11011001000111010100",

    "11011000110101101010",

    "11011000100100000010",

    "11011000010010011100",

    "11011000000000111001",

    "11010111101111010111",

    "11010111011101111000",

    "11010111001100011011",

    "11010110111011000000",

    "11010110101001100111",

    "11010110011000010000",

    "11010110000110111100",

    "11010101110101101001",

    "11010101100100011000",

    "11010101010011001010",

    "11010101000001111110",

    "11010100110000110011",

    "11010100011111101011",

    "11010100001110100101",

    "11010011111101100001",

    "11010011101100011111",

    "11010011011011011111",

    "11010011001010100001",

    "11010010111001100101",

    "11010010101000101011",

    "11010010010111110100",

    "11010010000110111110",

    "11010001110110001010",

    "11010001100101011000",

    "11010001010100101001",

    "11010001000011111011",

    "11010000110011001111",

    "11010000100010100101",

    "11010000010001111110",

    "11010000000001011000",

    "11001111110000110100",

    "11001111100000010010",

    "11001111001111110011",

    "11001110111111010101",

    "11001110101110111001",

    "11001110011110011111",

    "11001110001110000111",

    "11001101111101110001",

    "11001101101101011101",

    "11001101011101001011",

    "11001101001100111010",

    "11001100111100101100",

    "11001100101100100000",

    "11001100011100010101",

    "11001100001100001101",

    "11001011111100000110",

    "11001011101100000001",

    "11001011011011111110",

    "11001011001011111101",

    "11001010111011111110",

    "11001010101100000001",

    "11001010011100000110",

    "11001010001100001101",

    "11001001111100010101",

    "11001001101100011111",

    "11001001011100101100",

    "11001001001100111010",

    "11001000111101001001",

    "11001000101101011011",

    "11001000011101101111",

    "11001000001110000100",

    "11000111111110011100",

    "11000111101110110101",

    "11000111011111010000",

    "11000111001111101100",

    "11000111000000001011",

    "11000110110000101011",

    "11000110100001001101",

    "11000110010001110001",

    "11000110000010010111",

    "11000101110010111111",

    "11000101100011101000",

    "11000101010100010011",

    "11000101000101000000",

    "11000100110101101111",

    "11000100100110011111",

    "11000100010111010010",

    "11000100001000000110",

    "11000011111000111100",

    "11000011101001110011",

    "11000011011010101100",

    "11000011001011100111",

    "11000010111100100100",

    "11000010101101100011",

    "11000010011110100011",

    "11000010001111100101",

    "11000010000000101001",

    "11000001110001101110",

    "11000001100010110101",

    "11000001010011111110",

    "11000001000101001001",

    "11000000110110010101",

    "11000000100111100011",

    "11000000011000110011",

    "11000000001010000100",

    "10111111111011010111",

    "10111111101100101100",

    "10111111011110000011",

    "10111111001111011011",

    "10111111000000110100",

    "10111110110010010000",

    "10111110100011101101",

    "10111110010101001100",

    "10111110000110101100",

    "10111101111000001110",

    "10111101101001110010",

    "10111101011011011000",

    "10111101001100111111",

    "10111100111110100111",

    "10111100110000010010",

    "10111100100001111110",

    "10111100010011101011",

    "10111100000101011010",

    "10111011110111001011",

    "10111011101000111110",

    "10111011011010110010",

    "10111011001100100111",

    "10111010111110011111",

    "10111010110000011000",

    "10111010100010010010",

    "10111010010100001110",

    "10111010000110001100",

    "10111001111000001011",

    "10111001101010001100",

    "10111001011100001110",

    "10111001001110010010",

    "10111001000000011000",

    "10111000110010011111",

    "10111000100100100111",

    "10111000010110110010",

    "10111000001000111101",

    "10110111111011001011",

    "10110111101101011010",

    "10110111011111101010",

    "10110111010001111100",

    "10110111000100010000",

    "10110110110110100101",

    "10110110101000111011",

    "10110110011011010011",

    "10110110001101101101",

    "10110110000000001000",

    "10110101110010100101",

    "10110101100101000011",

    "10110101010111100011",

    "10110101001010000100",

    "10110100111100100110",

    "10110100101111001011",

    "10110100100001110000",

    "10110100010100010111",

    "10110100000111000000",

    "10110011111001101010",

    "10110011101100010110",

    "10110011011111000011",

    "10110011010001110010",

    "10110011000100100010",

    "10110010110111010011",

    "10110010101010000110",

    "10110010011100111011",

    "10110010001111110001",

    "10110010000010101000",

    "10110001110101100001",

    "10110001101000011011",

    "10110001011011010111",

    "10110001001110010100",

    "10110001000001010010",

    "10110000110100010010",

    "10110000100111010100",

    "10110000011010010111",

    "10110000001101011011",

    "10110000000000100001",

    "10101111110011101000",

    "10101111100110110000",

    "10101111011001111010",

    "10101111001101000110",

    "10101111000000010011",

    "10101110110011100001",

    "10101110100110110000",

    "10101110011010000001",

    "10101110001101010100",

    "10101110000000100111",

    "10101101110011111101",

    "10101101100111010011",

    "10101101011010101011",

    "10101101001110000100",

    "10101101000001011111",

    "10101100110100111011",

    "10101100101000011000",

    "10101100011011110111",

    "10101100001111010111",

    "10101100000010111001",

    "10101011110110011100",

    "10101011101010000000",

    "10101011011101100101",

    "10101011010001001100",

    "10101011000100110100",

    "10101010111000011110",

    "10101010101100001001",

    "10101010011111110101",

    "10101010010011100011",

    "10101010000111010001",

    "10101001111011000010",

    "10101001101110110011",

    "10101001100010100110",

    "10101001010110011010",

    "10101001001010010000",

    "10101000111110000111",

    "10101000110001111111",

    "10101000100101111000",

    "10101000011001110011",

    "10101000001101101111",

    "10101000000001101100",

    "10100111110101101011",

    "10100111101001101011",

    "10100111011101101100",

    "10100111010001101110",

    "10100111000101110010",

    "10100110111001110111",

    "10100110101101111101",

    "10100110100010000101",

    "10100110010110001110",

    "10100110001010011000",

    "10100101111110100011",

    "10100101110010110000",

    "10100101100110111101",

    "10100101011011001101",

    "10100101001111011101",

    "10100101000011101111",

    "10100100111000000010",

    "10100100101100010110",

    "10100100100000101011",

    "10100100010101000010",

    "10100100001001011001",

    "10100011111101110011",

    "10100011110010001101",

    "10100011100110101000",

    "10100011011011000101",

    "10100011001111100011",

    "10100011000100000010",

    "10100010111000100011",

    "10100010101101000100",

    "10100010100001100111",

    "10100010010110001011",

    "10100010001010110001",

    "10100001111111010111",

    "10100001110011111111",

    "10100001101000101000",

    "10100001011101010010",

    "10100001010001111101",

    "10100001000110101001",

    "10100000111011010111",

    "10100000110000000110",

    "10100000100100110110",

    "10100000011001100111",

    "10100000001110011001",

    "10100000000011001101",

    "10011111111000000010",

    "10011111101100110111",

    "10011111100001101110",

    "10011111010110100111",

    "10011111001011100000",

    "10011111000000011011",

    "10011110110101010110",

    "10011110101010010011",

    "10011110011111010001",

    "10011110010100010000",

    "10011110001001010001",

    "10011101111110010010",

    "10011101110011010101",

    "10011101101000011000",

    "10011101011101011101",

    "10011101010010100011",

    "10011101000111101010",

    "10011100111100110011",

    "10011100110001111100",

    "10011100100111000110",

    "10011100011100010010",

    "10011100010001011111",

    "10011100000110101101",

    "10011011111011111100",

    "10011011110001001100",

    "10011011100110011101",

    "10011011011011101111",

    "10011011010001000011",

    "10011011000110010111",

    "10011010111011101101",

    "10011010110001000100",

    "10011010100110011011",

    "10011010011011110100",

    "10011010010001001110",

    "10011010000110101001",

    "10011001111100000110",

    "10011001110001100011",

    "10011001100111000001",

    "10011001011100100001",

    "10011001010010000001",

    "10011001000111100011",

    "10011000111101000101",

    "10011000110010101001",

    "10011000101000001110",

    "10011000011101110100",

    "10011000010011011011",

    "10011000001001000011",

    "10010111111110101100",

    "10010111110100010110",

    "10010111101010000001",

    "10010111011111101101",

    "10010111010101011011",

    "10010111001011001001",

    "10010111000000111000",

    "10010110110110101001",

    "10010110101100011010",

    "10010110100010001101",

    "10010110011000000000",

    "10010110001101110101",

    "10010110000011101010",

    "10010101111001100001",

    "10010101101111011001",

    "10010101100101010001",

    "10010101011011001011",

    "10010101010001000110",

    "10010101000111000001",

    "10010100111100111110",

    "10010100110010111100",

    "10010100101000111011",

    "10010100011110111011",

    "10010100010100111011",

    "10010100001010111101",

    "10010100000001000000",

    "10010011110111000100",

    "10010011101101001001",

    "10010011100011001110",

    "10010011011001010101",

    "10010011001111011101",

    "10010011000101100110",

    "10010010111011110000",

    "10010010110001111011",

    "10010010101000000110",

    "10010010011110010011",

    "10010010010100100001",

    "10010010001010110000",

    "10010010000000111111",

    "10010001110111010000",

    "10010001101101100010",

    "10010001100011110100",

    "10010001011010001000",

    "10010001010000011100",

    "10010001000110110010",

    "10010000111101001000",

    "10010000110011100000",

    "10010000101001111000",

    "10010000100000010010",

    "10010000010110101100",

    "10010000001101000111",

    "10010000000011100011",

    "10001111111010000001",

    "10001111110000011111",

    "10001111100110111110",

    "10001111011101011110",

    "10001111010011111111",

    "10001111001010100001",

    "10001111000001000011",

    "10001110110111100111",

    "10001110101110001100",

    "10001110100100110010",

    "10001110011011011000",

    "10001110010010000000",

    "10001110001000101000",

    "10001101111111010001",

    "10001101110101111100",

    "10001101101100100111",

    "10001101100011010011",

    "10001101011010000000",

    "10001101010000101110",

    "10001101000111011101",

    "10001100111110001101",

    "10001100110100111101",

    "10001100101011101111",

    "10001100100010100001",

    "10001100011001010101",

    "10001100010000001001",

    "10001100000110111110",

    "10001011111101110100",

    "10001011110100101011",

    "10001011101011100011",

    "10001011100010011100",

    "10001011011001010110",

    "10001011010000010000",

    "10001011000111001100",

    "10001010111110001000",

    "10001010110101000101",

    "10001010101100000100",

    "10001010100011000011",

    "10001010011010000010",

    "10001010010001000011",

    "10001010001000000101",

    "10001001111111000111",

    "10001001110110001011",

    "10001001101101001111",

    "10001001100100010100",

    "10001001011011011010",

    "10001001010010100001",

    "10001001001001101000",

    "10001001000000110001",

    "10001000110111111010",

    "10001000101111000101",

    "10001000100110010000",

    "10001000011101011100",

    "10001000010100101001",

    "10001000001011110110",

    "10001000000011000101",

    "10000111111010010100",

    "10000111110001100100",

    "10000111101000110110",

    "10000111100000000111",

    "10000111010111011010",

    "10000111001110101110",

    "10000111000110000010",

    "10000110111101010111",

    "10000110110100101110",

    "10000110101100000101",

    "10000110100011011100",

    "10000110011010110101",

    "10000110010010001110",

    "10000110001001101001",

    "10000110000001000100",

    "10000101111000011111",

    "10000101101111111100",

    "10000101100111011010",

    "10000101011110111000",

    "10000101010110010111",

    "10000101001101110111",

    "10000101000101011000",

    "10000100111100111010",

    "10000100110100011100",

    "10000100101011111111",

    "10000100100011100011",

    "10000100011011001000",

    "10000100010010101110",

    "10000100001010010100",

    "10000100000001111011",

    "10000011111001100011",

    "10000011110001001100",

    "10000011101000110110",

    "10000011100000100000",

    "10000011011000001011",

    "10000011001111110111",

    "10000011000111100100",

    "10000010111111010010",

    "10000010110111000000",

    "10000010101110101111",

    "10000010100110011111",

    "10000010011110010000",

    "10000010010110000001",

    "10000010001101110100",

    "10000010000101100111",

    "10000001111101011011",

    "10000001110101001111",

    "10000001101101000100",

    "10000001100100111011",

    "10000001011100110001",

    "10000001010100101001",

    "10000001001100100010",

    "10000001000100011011",

    "10000000111100010101",

    "10000000110100001111",

    "10000000101100001011",

    "10000000100100000111",

    "10000000011100000100",

    "10000000010100000010",

    "10000000001100000000",

    "10000000000100000000"
	);
	
begin

main_proc: process(rom_enable)

begin


if(rom_enable = '1') then

data_out <= mem(to_integer(unsigned(address)));

end if;

end process;

end architecture;