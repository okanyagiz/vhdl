library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.all;
use IEEE.NUMERIC_STD.ALL;

entity my_rom_dp is 
generic(

addr_len: natural := 10;
data_len: natural := 20
);
port(
rom_enable: in std_logic;
address: in std_logic_vector((addr_len -1) downto 0);
data_out: out std_logic_vector((data_len -1) downto 0)
);
end entity;


architecture arch of my_rom_dp is

type rom_type is array (0 to (2**(addr_len) -1)) of std_logic_vector((data_len -1) downto 0);

constant mem: rom_type := 
	(
	"11111111100000000001",

    "11111110100000001101",

    "11111101100000100101",

    "11111100100001001001",

    "11111011100001111000",

    "11111010100010110100",

    "11111001100011111011",

    "11111000100101001110",

    "11110111100110101100",

    "11110110101000010110",

    "11110101101010001100",

    "11110100101100001101",

    "11110011101110011010",

    "11110010110000110010",

    "11110001110011010110",

    "11110000110110000100",

    "11101111111000111111",

    "11101110111100000100",

    "11101101111111010101",

    "11101101000010110000",

    "11101100000110010111",

    "11101011001010001001",

    "11101010001110000110",

    "11101001010010001110",

    "11101000010110100001",

    "11100111011010111111",

    "11100110011111101000",

    "11100101100100011100",

    "11100100101001011010",

    "11100011101110100011",

    "11100010110011110111",

    "11100001111001010110",

    "11100000111110111111",

    "11100000000100110011",

    "11011111001010110001",

    "11011110010000111010",

    "11011101010111001101",

    "11011100011101101011",

    "11011011100100010011",

    "11011010101011000110",

    "11011001110010000011",

    "11011000111001001010",

    "11011000000000011011",

    "11010111000111110110",

    "11010110001111011100",

    "11010101010111001100",

    "11010100011111000110",

    "11010011100111001010",

    "11010010101111011000",

    "11010001110111110000",

    "11010001000000010001",

    "11010000001000111101",

    "11001111010001110011",

    "11001110011010110010",

    "11001101100011111011",

    "11001100101101001110",

    "11001011110110101011",

    "11001011000000010001",

    "11001010001010000001",

    "11001001010011111011",

    "11001000011101111110",

    "11000111101000001011",

    "11000110110010100001",

    "11000101111101000001",

    "11000101000111101010",

    "11000100010010011101",

    "11000011011101011000",

    "11000010101000011110",

    "11000001110011101100",

    "11000000111111000100",

    "11000000001010100101",

    "10111111010110001111",

    "10111110100010000011",

    "10111101101101111111",

    "10111100111010000101",

    "10111100000110010011",

    "10111011010010101011",

    "10111010011111001100",

    "10111001101011110101",

    "10111000111000101000",

    "10111000000101100011",

    "10110111010010101000",

    "10110110011111110101",

    "10110101101101001011",

    "10110100111010101010",

    "10110100001000010001",

    "10110011010110000001",

    "10110010100011111010",

    "10110001110001111100",

    "10110001000000000110",

    "10110000001110011000",

    "10101111011100110100",

    "10101110101011010111",

    "10101101111010000100",

    "10101101001000111000",

    "10101100010111110110",

    "10101011100110111011",

    "10101010110110001001",

    "10101010000101011111",

    "10101001010100111110",

    "10101000100100100101",

    "10100111110100010100",

    "10100111000100001011",

    "10100110010100001011",

    "10100101100100010010",

    "10100100110100100010",

    "10100100000100111010",

    "10100011010101011010",

    "10100010100110000010",

    "10100001110110110010",

    "10100001000111101010",

    "10100000011000101011",

    "10011111101001110010",

    "10011110111011000010",

    "10011110001100011010",

    "10011101011101111010",

    "10011100101111100001",

    "10011100000001010000",

    "10011011010011000111",

    "10011010100101000110",

    "10011001110111001101",

    "10011001001001011011",

    "10011000011011110001",

    "10010111101110001110",

    "10010111000000110011",

    "10010110010011100000",

    "10010101100110010100",

    "10010100111001010000",

    "10010100001100010011",

    "10010011011111011110",

    "10010010110010110000",

    "10010010000110001010",

    "10010001011001101011",

    "10010000101101010011",

    "10010000000001000011",

    "10001111010100111010",

    "10001110101000111000",

    "10001101111100111110",

    "10001101010001001011",

    "10001100100101011111",

    "10001011111001111010",

    "10001011001110011100",

    "10001010100011000110",

    "10001001110111110111",

    "10001001001100101111",

    "10001000100001101110",

    "10000111110110110100",

    "10000111001100000001",

    "10000110100001010101",

    "10000101110110110000",

    "10000101001100010010",

    "10000100100001111011",

    "10000011110111101010",

    "10000011001101100001",

    "10000010100011011111",

    "10000001111001100011",

    "10000001001111101110",

    "10000000100110000000",

    "01111111111100011001",

    "01111111010010111001",

    "01111110101001011111",

    "01111110000000001100",

    "01111101010110111111",

    "01111100101101111010",

    "01111100000100111011",

    "01111011011100000010",

    "01111010110011010000",

    "01111010001010100101",

    "01111001100010000000",

    "01111000111001100010",

    "01111000010001001010",

    "01110111101000111001",

    "01110111000000101110",

    "01110110011000101010",

    "01110101110000101100",

    "01110101001000110100",

    "01110100100001000011",

    "01110011111001011000",

    "01110011010001110100",

    "01110010101010010110",

    "01110010000010111110",

    "01110001011011101100",

    "01110000110100100001",

    "01110000001101011100",

    "01101111100110011101",

    "01101110111111100100",

    "01101110011000110001",

    "01101101110010000101",

    "01101101001011011111",

    "01101100100100111110",

    "01101011111110100100",

    "01101011011000010000",

    "01101010110010000010",

    "01101010001011111010",

    "01101001100101111000",

    "01101000111111111100",

    "01101000011010000110",

    "01100111110100010110",

    "01100111001110101100",

    "01100110101001001000",

    "01100110000011101001",

    "01100101011110010001",

    "01100100111000111110",

    "01100100010011110001",

    "01100011101110101010",

    "01100011001001101001",

    "01100010100100101110",

    "01100001111111111000",

    "01100001011011001000",

    "01100000110110011110",

    "01100000010001111001",

    "01011111101101011011",

    "01011111001001000001",

    "01011110100100101110",

    "01011110000000100000",

    "01011101011100011000",

    "01011100111000010101",

    "01011100010100011000",

    "01011011110000100000",

    "01011011001100101110",

    "01011010101001000010",

    "01011010000101011010",

    "01011001100001111001",

    "01011000111110011101",

    "01011000011011000110",

    "01010111110111110101",

    "01010111010100101001",

    "01010110110001100011",

    "01010110001110100010",

    "01010101101011100110",

    "01010101001000110000",

    "01010100100101111111",

    "01010100000011010011",

    "01010011100000101101",

    "01010010111110001100",

    "01010010011011110000",

    "01010001111001011001",

    "01010001010111001000",

    "01010000110100111100",

    "01010000010010110101",

    "01001111110000110011",

    "01001111001110110110",

    "01001110101100111111",

    "01001110001011001100",

    "01001101101001011111",

    "01001101000111110111",

    "01001100100110010100",

    "01001100000100110110",

    "01001011100011011101",

    "01001011000010001001",

    "01001010100000111010",

    "01001001111111110000",

    "01001001011110101011",

    "01001000111101101011",

    "01001000011100110000",

    "01000111111011111010",

    "01000111011011001001",

    "01000110111010011101",

    "01000110011001110101",

    "01000101111001010011",

    "01000101011000110101",

    "01000100111000011100",

    "01000100011000001000",

    "01000011110111111001",

    "01000011010111101111",

    "01000010110111101001",

    "01000010010111101001",

    "01000001110111101101",

    "01000001010111110101",

    "01000000111000000011",

    "01000000011000010101",

    "00111111111000101100",

    "00111111011001001000",

    "00111110111001101000",

    "00111110011010001101",

    "00111101111010110110",

    "00111101011011100100",

    "00111100111100010111",

    "00111100011101001110",

    "00111011111110001010",

    "00111011011111001011",

    "00111011000000010000",

    "00111010100001011010",

    "00111010000010101000",

    "00111001100011111010",

    "00111001000101010010",

    "00111000100110101101",

    "00111000001000001101",

    "00110111101001110010",

    "00110111001011011011",

    "00110110101101001001",

    "00110110001110111010",

    "00110101110000110001",

    "00110101010010101011",

    "00110100110100101010",

    "00110100010110101110",

    "00110011111000110110",

    "00110011011011000010",

    "00110010111101010010",

    "00110010011111100111",

    "00110010000010000000",

    "00110001100100011101",

    "00110001000110111111",

    "00110000101001100101",

    "00110000001100001111",

    "00101111101110111101",

    "00101111010001110000",

    "00101110110100100111",

    "00101110010111100010",

    "00101101111010100001",

    "00101101011101100100",

    "00101101000000101100",

    "00101100100011110111",

    "00101100000111000111",

    "00101011101010011011",

    "00101011001101110011",

    "00101010110001001111",

    "00101010010100110000",

    "00101001111000010100",

    "00101001011011111100",

    "00101000111111101001",

    "00101000100011011001",

    "00101000000111001101",

    "00100111101011000110",

    "00100111001111000010",

    "00100110110011000011",

    "00100110010111000111",

    "00100101111011010000",

    "00100101011111011100",

    "00100101000011101100",

    "00100100101000000001",

    "00100100001100011001",

    "00100011110000110101",

    "00100011010101010101",

    "00100010111001111001",

    "00100010011110100000",

    "00100010000011001100",

    "00100001100111111100",

    "00100001001100101111",

    "00100000110001100110",

    "00100000010110100001",

    "00011111111011100000",

    "00011111100000100010",

    "00011111000101101000",

    "00011110101010110010",

    "00011110010000000000",

    "00011101110101010010",

    "00011101011010100111",

    "00011101000000000000",

    "00011100100101011101",

    "00011100001010111110",

    "00011011110000100010",

    "00011011010110001010",

    "00011010111011110101",

    "00011010100001100100",

    "00011010000111010111",

    "00011001101101001110",

    "00011001010011001000",

    "00011000111001000110",

    "00011000011111000111",

    "00011000000101001100",

    "00010111101011010101",

    "00010111010001100001",

    "00010110110111110001",

    "00010110011110000100",

    "00010110000100011011",

    "00010101101010110101",

    "00010101010001010011",

    "00010100110111110100",

    "00010100011110011001",

    "00010100000101000010",

    "00010011101011101110",

    "00010011010010011101",

    "00010010111001010000",

    "00010010100000000110",

    "00010010000111000000",

    "00010001101101111101",

    "00010001010100111110",

    "00010000111100000010",

    "00010000100011001001",

    "00010000001010010100",

    "00001111110001100010",

    "00001111011000110100",

    "00001111000000001001",

    "00001110100111100010",

    "00001110001110111101",

    "00001101110110011100",

    "00001101011101111111",

    "00001101000101100100",

    "00001100101101001110",

    "00001100010100111010",

    "00001011111100101010",

    "00001011100100011100",

    "00001011001100010011",

    "00001010110100001100",

    "00001010011100001001",

    "00001010000100001001",

    "00001001101100001100",

    "00001001010100010011",

    "00001000111100011100",

    "00001000100100101001",

    "00001000001100111001",

    "00000111110101001101",

    "00000111011101100011",

    "00000111000101111101",

    "00000110101110011001",

    "00000110010110111001",

    "00000101111111011101",

    "00000101101000000011",

    "00000101010000101100",

    "00000100111001011001",

    "00000100100010001000",

    "00000100001010111011",

    "00000011110011110001",

    "00000011011100101010",

    "00000011000101100110",

    "00000010101110100101",

    "00000010010111100111",

    "00000010000000101101",

    "00000001101001110101",

    "00000001010011000000",

    "00000000111100001110",

    "00000000100101100000",

    "00000000001110110100",

    "11111111110000011000",

    "11111111000011001100",

    "11111110010110000111",

    "11111101101001001000",

    "11111100111100001111",

    "11111100001111011011",

    "11111011100010101110",

    "11111010110110000110",

    "11111010001001100100",

    "11111001011101001000",

    "11111000110000110010",

    "11111000000100100010",

    "11110111011000011000",

    "11110110101100010011",

    "11110110000000010100",

    "11110101010100011011",

    "11110100101000101000",

    "11110011111100111010",

    "11110011010001010011",

    "11110010100101110001",

    "11110001111010010100",

    "11110001001110111101",

    "11110000100011101100",

    "11101111111000100001",

    "11101111001101011011",

    "11101110100010011011",

    "11101101110111100000",

    "11101101001100101011",

    "11101100100001111100",

    "11101011110111010010",

    "11101011001100101101",

    "11101010100010001111",

    "11101001110111110101",

    "11101001001101100001",

    "11101000100011010011",

    "11100111111001001010",

    "11100111001111000111",

    "11100110100101001001",

    "11100101111011010000",

    "11100101010001011101",

    "11100100100111101111",

    "11100011111110000111",

    "11100011010100100011",

    "11100010101011000110",

    "11100010000001101101",

    "11100001011000011010",

    "11100000101111001100",

    "11100000000110000100",

    "11011111011101000001",

    "11011110110100000011",

    "11011110001011001010",

    "11011101100010010111",

    "11011100111001101000",

    "11011100010000111111",

    "11011011101000011011",

    "11011010111111111101",

    "11011010010111100011",

    "11011001101111001111",

    "11011001000111000000",

    "11011000011110110110",

    "11010111110110110001",

    "11010111001110110001",

    "11010110100110110110",

    "11010101111111000000",

    "11010101010111001111",

    "11010100101111100100",

    "11010100000111111101",

    "11010011100000011100",

    "11010010111000111111",

    "11010010010001100111",

    "11010001101010010101",

    "11010001000011000111",

    "11010000011011111110",

    "11001111110100111011",

    "11001111001101111100",

    "11001110100111000010",

    "11001110000000001101",

    "11001101011001011101",

    "11001100110010110001",

    "11001100001100001011",

    "11001011100101101001",

    "11001010111111001101",

    "11001010011000110101",

    "11001001110010100001",

    "11001001001100010011",

    "11001000100110001010",

    "11001000000000000101",

    "11000111011010000101",

    "11000110110100001010",

    "11000110001110010011",

    "11000101101000100001",

    "11000101000010110100",

    "11000100011101001100",

    "11000011110111101000",

    "11000011010010001001",

    "11000010101100101111",

    "11000010000111011001",

    "11000001100010001000",

    "11000000111100111011",

    "11000000010111110100",

    "10111111110010110000",

    "10111111001101110010",

    "10111110101000111000",

    "10111110000100000010",

    "10111101011111010001",

    "10111100111010100101",

    "10111100010101111101",

    "10111011110001011001",

    "10111011001100111011",

    "10111010101000100000",

    "10111010000100001010",

    "10111001011111111001",

    "10111000111011101100",

    "10111000010111100011",

    "10110111110011011111",

    "10110111001111100000",

    "10110110101011100101",

    "10110110000111101110",

    "10110101100011111011",

    "10110101000000001101",

    "10110100011100100100",

    "10110011111000111110",

    "10110011010101011101",

    "10110010110010000001",

    "10110010001110101000",

    "10110001101011010100",

    "10110001001000000101",

    "10110000100100111001",

    "10110000000001110010",

    "10101111011110101111",

    "10101110111011110001",

    "10101110011000110111",

    "10101101110110000001",

    "10101101010011001111",

    "10101100110000100001",

    "10101100001101111000",

    "10101011101011010010",

    "10101011001000110001",

    "10101010100110010101",

    "10101010000011111100",

    "10101001100001100111",

    "10101000111111010111",

    "10101000011101001011",

    "10100111111011000011",

    "10100111011000111111",

    "10100110110110111111",

    "10100110010101000011",

    "10100101110011001011",

    "10100101010001010111",

    "10100100101111101000",

    "10100100001101111100",

    "10100011101100010101",

    "10100011001010110001",

    "10100010101001010010",

    "10100010000111110110",

    "10100001100110011111",

    "10100001000101001011",

    "10100000100011111100",

    "10100000000010110000",

    "10011111100001101001",

    "10011111000000100101",

    "10011110011111100110",

    "10011101111110101010",

    "10011101011101110010",

    "10011100111100111110",

    "10011100011100001110",

    "10011011111011100010",

    "10011011011010111010",

    "10011010111010010110",

    "10011010011001110101",

    "10011001111001011001",

    "10011001011001000000",

    "10011000111000101011",

    "10011000011000011010",

    "10010111111000001100",

    "10010111011000000011",

    "10010110110111111101",

    "10010110010111111011",

    "10010101110111111101",

    "10010101011000000011",

    "10010100111000001100",

    "10010100011000011010",

    "10010011111000101011",

    "10010011011000111111",

    "10010010111001011000",

    "10010010011001110100",

    "10010001111010010011",

    "10010001011010110111",

    "10010000111011011110",

    "10010000011100001001",

    "10001111111100111000",

    "10001111011101101010",

    "10001110111110100000",

    "10001110011111011001",

    "10001110000000010110",

    "10001101100001010111",

    "10001101000010011011",

    "10001100100011100011",

    "10001100000100101111",

    "10001011100101111110",

    "10001011000111010001",

    "10001010101000100111",

    "10001010001010000001",

    "10001001101011011110",

    "10001001001100111111",

    "10001000101110100100",

    "10001000010000001100",

    "10000111110001111000",

    "10000111010011100111",

    "10000110110101011001",

    "10000110010111001111",

    "10000101111001001001",

    "10000101011011000110",

    "10000100111101000111",

    "10000100011111001011",

    "10000100000001010010",

    "10000011100011011101",

    "10000011000101101011",

    "10000010100111111101",

    "10000010001010010010",

    "10000001101100101011",

    "10000001001111000111",

    "10000000110001100110",

    "10000000010100001001",

    "01111111110110101111",

    "01111111011001011001",

    "01111110111100000110",

    "01111110011110110110",

    "01111110000001101001",

    "01111101100100100000",

    "01111101000111011011",

    "01111100101010011000",

    "01111100001101011001",

    "01111011110000011101",

    "01111011010011100101",

    "01111010110110110000",

    "01111010011001111110",

    "01111001111101001111",

    "01111001100000100100",

    "01111001000011111100",

    "01111000100111010111",

    "01111000001010110101",

    "01110111101110010111",

    "01110111010001111100",

    "01110110110101100100",

    "01110110011001001111",

    "01110101111100111110",

    "01110101100000110000",

    "01110101000100100101",

    "01110100101000011101",

    "01110100001100011000",

    "01110011110000010110",

    "01110011010100011000",

    "01110010111000011101",

    "01110010011100100101",

    "01110010000000110000",

    "01110001100100111110",

    "01110001001001001111",

    "01110000101101100100",

    "01110000010001111011",

    "01101111110110010110",

    "01101111011010110100",

    "01101110111111010101",

    "01101110100011111001",

    "01101110001000100000",

    "01101101101101001010",

    "01101101010001110111",

    "01101100110110100111",

    "01101100011011011010",

    "01101100000000010001",

    "01101011100101001010",

    "01101011001010000110",

    "01101010101111000110",

    "01101010010100001000",

    "01101001111001001101",

    "01101001011110010110",

    "01101001000011100001",

    "01101000101000101111",

    "01101000001110000001",

    "01100111110011010101",

    "01100111011000101100",

    "01100110111110000111",

    "01100110100011100100",

    "01100110001001000100",

    "01100101101110100111",

    "01100101010100001101",

    "01100100111001110110",

    "01100100011111100010",

    "01100100000101010000",

    "01100011101011000010",

    "01100011010000110110",

    "01100010110110101110",

    "01100010011100101000",

    "01100010000010100101",

    "01100001101000100101",

    "01100001001110101000",

    "01100000110100101110",

    "01100000011010110111",

    "01100000000001000010",

    "01011111100111010000",

    "01011111001101100001",

    "01011110110011110101",

    "01011110011010001100",

    "01011110000000100110",

    "01011101100111000010",

    "01011101001101100001",

    "01011100110100000011",

    "01011100011010101000",

    "01011100000001001111",

    "01011011100111111010",

    "01011011001110100111",

    "01011010110101010110",

    "01011010011100001001",

    "01011010000010111110",

    "01011001101001110110",

    "01011001010000110001",

    "01011000110111101111",

    "01011000011110101111",

    "01011000000101110010",

    "01010111101100111000",

    "01010111010100000000",

    "01010110111011001011",

    "01010110100010011001",

    "01010110001001101001",

    "01010101110000111100",

    "01010101011000010010",

    "01010100111111101011",

    "01010100100111000110",

    "01010100001110100011",

    "01010011110110000100",

    "01010011011101100111",

    "01010011000101001101",

    "01010010101100110101",

    "01010010010100100000",

    "01010001111100001110",

    "01010001100011111110",

    "01010001001011110001",

    "01010000110011100110",

    "01010000011011011110",

    "01010000000011011001",

    "01001111101011010110",

    "01001111010011010110",

    "01001110111011011000",

    "01001110100011011101",

    "01001110001011100100",

    "01001101110011101110",

    "01001101011011111011",

    "01001101000100001010",

    "01001100101100011100",

    "01001100010100110000",

    "01001011111101000110",

    "01001011100101100000",

    "01001011001101111011",

    "01001010110110011010",

    "01001010011110111010",

    "01001010000111011110",

    "01001001110000000100",

    "01001001011000101100",

    "01001001000001010111",

    "01001000101010000100",

    "01001000010010110011",

    "01000111111011100110",

    "01000111100100011010",

    "01000111001101010001",

    "01000110110110001011",

    "01000110011111000111",

    "01000110001000000101",

    "01000101110001000110",

    "01000101011010001001",

    "01000101000011001111",

    "01000100101100010111",

    "01000100010101100010",

    "01000011111110101111",

    "01000011100111111110",

    "01000011010001010000",

    "01000010111010100100",

    "01000010100011111010",

    "01000010001101010011",

    "01000001110110101110",

    "01000001100000001100",

    "01000001001001101100",

    "01000000110011001110",

    "01000000011100110011",

    "01000000000110011010",

    "00111111110000000100",

    "00111111011001101111",

    "00111111000011011101",

    "00111110101101001110",

    "00111110010111000001",

    "00111110000000110110",

    "00111101101010101101",

    "00111101010100100111",

    "00111100111110100011",

    "00111100101000100001",

    "00111100010010100010",

    "00111011111100100100",

    "00111011100110101010",

    "00111011010000110001",

    "00111010111010111011",

    "00111010100101000111",

    "00111010001111010101",

    "00111001111001100110",

    "00111001100011111000",

    "00111001001110001101",

    "00111000111000100101",

    "00111000100010111110",

    "00111000001101011010",

    "00110111110111111000",

    "00110111100010011000",

    "00110111001100111010",

    "00110110110111011111",

    "00110110100010000110",

    "00110110001100101111",

    "00110101110111011010",

    "00110101100010001000",

    "00110101001100110111",

    "00110100110111101001",

    "00110100100010011101",

    "00110100001101010011",

    "00110011111000001100",

    "00110011100011000110",

    "00110011001110000011",

    "00110010111001000010",

    "00110010100100000011",

    "00110010001111000110",

    "00110001111010001011",

    "00110001100101010011",

    "00110001010000011100",

    "00110000111011101000",

    "00110000100110110110",

    "00110000010010000110",

    "00101111111101011000",

    "00101111101000101100",

    "00101111010100000011",

    "00101110111111011011",

    "00101110101010110110",

    "00101110010110010010",

    "00101110000001110001",

    "00101101101101010010",

    "00101101011000110101",

    "00101101000100011010",

    "00101100110000000001",

    "00101100011011101010",

    "00101100000111010101",

    "00101011110011000010",

    "00101011011110110010",

    "00101011001010100011",

    "00101010110110010110",

    "00101010100010001100",

    "00101010001110000011",

    "00101001111001111101",

    "00101001100101111000",

    "00101001010001110110",

    "00101000111101110110",

    "00101000101001110111",

    "00101000010101111011",

    "00101000000010000000",

    "00100111101110001000",

    "00100111011010010010",

    "00100111000110011101",

    "00100110110010101011",

    "00100110011110111011",

    "00100110001011001100",

    "00100101110111100000",

    "00100101100011110110",

    "00100101010000001101",

    "00100100111100100111",

    "00100100101001000010",

    "00100100010101100000",

    "00100100000001111111",

    "00100011101110100000",

    "00100011011011000100",

    "00100011000111101001",

    "00100010110100010000",

    "00100010100000111001",

    "00100010001101100100",

    "00100001111010010001",

    "00100001100111000000",

    "00100001010011110001",

    "00100001000000100100",

    "00100000101101011000",

    "00100000011010001111",

    "00100000000111000111",

    "00011111110100000010",

    "00011111100000111110",

    "00011111001101111100",

    "00011110111010111100",

    "00011110100111111110",

    "00011110010101000010",

    "00011110000010000111",

    "00011101101111001111",

    "00011101011100011000",

    "00011101001001100100",

    "00011100110110110001",

    "00011100100100000000",

    "00011100010001010001",

    "00011011111110100011",

    "00011011101011111000",

    "00011011011001001110",

    "00011011000110100111",

    "00011010110100000001",

    "00011010100001011101",

    "00011010001110111010",

    "00011001111100011010",

    "00011001101001111011",

    "00011001010111011110",

    "00011001000101000011",

    "00011000110010101010",

    "00011000100000010011",

    "00011000001101111101",

    "00010111111011101001",

    "00010111101001010111",

    "00010111010111000111",

    "00010111000100111001",

    "00010110110010101100",

    "00010110100000100001",

    "00010110001110011000",

    "00010101111100010001",

    "00010101101010001011",

    "00010101011000001000",

    "00010101000110000110",

    "00010100110100000101",

    "00010100100010000111",

    "00010100010000001010",

    "00010011111110001111",

    "00010011101100010110",

    "00010011011010011110",

    "00010011001000101000",

    "00010010110110110100",

    "00010010100101000010",

    "00010010010011010001",

    "00010010000001100010",

    "00010001101111110101",

    "00010001011110001010",

    "00010001001100100000",

    "00010000111010111000",

    "00010000101001010010",

    "00010000010111101101",

    "00010000000110001010",

    "00001111110100101001",

    "00001111100011001001",

    "00001111010001101100",

    "00001111000000001111",

    "00001110101110110101",

    "00001110011101011100",

    "00001110001100000101",

    "00001101111010101111",

    "00001101101001011100",

    "00001101011000001010",

    "00001101000110111001",

    "00001100110101101010",

    "00001100100100011101",

    "00001100010011010010",

    "00001100000010001000",

    "00001011110000111111",

    "00001011011111111001",

    "00001011001110110100",

    "00001010111101110001",

    "00001010101100101111",

    "00001010011011101111",

    "00001010001010110001",

    "00001001111001110100",

    "00001001101000111001",

    "00001001010111111111",

    "00001001000111000111",

    "00001000110110010001",

    "00001000100101011100",

    "00001000010100101001",

    "00001000000011110111",

    "00000111110011000111",

    "00000111100010011001",

    "00000111010001101100",

    "00000111000001000001",

    "00000110110000010111",

    "00000110011111101111",

    "00000110001111001001",

    "00000101111110100100",

    "00000101101110000001",

    "00000101011101011111",

    "00000101001100111111",

    "00000100111100100000",

    "00000100101100000011",

    "00000100011011101000",

    "00000100001011001110",

    "00000011111010110110",

    "00000011101010011111",

    "00000011011010001001",

    "00000011001001110110",

    "00000010111001100011",

    "00000010101001010011",

    "00000010011001000100",

    "00000010001000110110",

    "00000001111000101010",

    "00000001101000011111",

    "00000001011000010110",

    "00000001001000001111",

    "00000000111000001001",

    "00000000101000000100",

    "00000000011000000001",

    "00000000001000000000"

	);
	
begin

main_proc: process(rom_enable)

begin


if(rom_enable = '1') then

data_out <= mem(to_integer(unsigned(address)));

end if;

end process;

end architecture;